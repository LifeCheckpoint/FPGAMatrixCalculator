`timescale 1ns / 1ps

module transform_3x3x4x4_8x10 (
    input  logic [15:0] tile  [0:2][0:2][0:3][0:3],
    output logic [15:0] image [0:7][0:9]
);

// In this module, input will be stick and clip invalid areas, not div.

always_comb begin
    image = '{
        tile[0][0][0][0], tile[0][0][0][1], tile[0][0][0][2], tile[0][0][0][3], tile[0][1][0][0], tile[0][1][0][1], tile[0][1][0][2], tile[0][1][0][3], tile[0][2][0][0], tile[0][2][0][1],
        tile[0][0][1][0], tile[0][0][1][1], tile[0][0][1][2], tile[0][0][1][3], tile[0][1][1][0], tile[0][1][1][1], tile[0][1][1][2], tile[0][1][1][3], tile[0][2][1][0], tile[0][2][1][1],
        tile[0][0][2][0], tile[0][0][2][1], tile[0][0][2][2], tile[0][0][2][3], tile[0][1][2][0], tile[0][1][2][1], tile[0][1][2][2], tile[0][1][2][3], tile[0][2][2][0], tile[0][2][2][1],
        tile[0][0][3][0], tile[0][0][3][1], tile[0][0][3][2], tile[0][0][3][3], tile[0][1][3][0], tile[0][1][3][1], tile[0][1][3][2], tile[0][1][3][3], tile[0][2][3][0], tile[0][2][3][1],
        tile[1][0][0][0], tile[1][0][0][1], tile[1][0][0][2], tile[1][0][0][3], tile[1][1][0][0], tile[1][1][0][1], tile[1][1][0][2], tile[1][1][0][3], tile[1][2][0][0], tile[1][2][0][1],
        tile[1][0][1][0], tile[1][0][1][1], tile[1][0][1][2], tile[1][0][1][3], tile[1][1][1][0], tile[1][1][1][1], tile[1][1][1][2], tile[1][1][1][3], tile[1][2][1][0], tile[1][2][1][1],
        tile[1][0][2][0], tile[1][0][2][1], tile[1][0][2][2], tile[1][0][2][3], tile[1][1][2][0], tile[1][1][2][1], tile[1][1][2][2], tile[1][1][2][3], tile[1][2][2][0], tile[1][2][2][1],
        tile[1][0][3][0], tile[1][0][3][1], tile[1][0][3][2], tile[1][0][3][3], tile[1][1][3][0], tile[1][1][3][1], tile[1][1][3][2], tile[1][1][3][3], tile[1][2][3][0], tile[1][2][3][1]
    };
end

endmodule
